// SYNTHESIZABLE ADDER FOR N BIT SIGNED MAGNITUDE WITH F BITS OF FRACTION
// CREATED BY MEHDI SAFAEE, WINTER 2018-2019
`include "config.svh"
module sigma8
//##############################################################################################
//##############################################################################################
// PARAMETERs-----------------------------------------------------------------------------------
// INPUT AND OUTPUTS----------------------------------------------------------------------------
    (
    input logic [`N-1:0] a0, a1, a2, a3, a4, a5, a6, a7,
    output logic [`N-1:0] c
    );
// MODULES INSTANTIATIONS-----------------------------------------------------------------------
    logic [`N-1:0] temp [0:1];
    logic [`N-1:0] result;

	sigma4 sigma4_0 
    (
		.a0(a0), .a1(a1), .a2(a2), .a3(a3), 
		.c(temp[0])
	);
    sigma4 sigma4_1
    (
		.a0(a4), .a1(a5), .a2(a6), .a3(a7),
		.c(temp[1])
	);
	adder adder0
    (
		.a(temp[0]), 
		.b(temp[1]), 
		.c(result)
	);
// VARIABLES -----------------------------------------------------------------------------------
    assign c = result;
// INITIALIZATIONS------------------------------------------------------------------------------
// MAIN-----------------------------------------------------------------------------------------
//##############################################################################################
//##############################################################################################
endmodule