// SYNTHESIZABLE MULTIPLIER FOR N BIT SIGNED MAGNITUDE WITH F BITS OF FRACTION
// CREATED BY MEHDI SAFAEE, WINTER 2018-2019
`include "config.svh"
module mask 
//##############################################################################################
//##############################################################################################
// PARAMETERs-----------------------------------------------------------------------------------
	#(
	parameter R = 3,
	parameter C = 4
	)
// INPUT AND OUTPUTS----------------------------------------------------------------------------
	(
	 input logic		[`nStates-1:0]	a,
	 					[`N-1:0] 		b[0:R-1][0:C-1],
	 output	logic		[`N-1:0]		c[0:R-1][0:C-1]
	 );
// VARIABLES -----------------------------------------------------------------------------------
// MODULES INSTANTIATIONS-----------------------------------------------------------------------
genvar i, j;
generate
	for (i=0; i<R; i=i+1) begin : loop_on_rows
	    for (j=0; j<C; j=j+1) begin : loop_on_columns
            assign c[i][j] = {`N{a[i]}} & b[i][j];
	end
	end
endgenerate
// INITIALIZATIONS------------------------------------------------------------------------------	
// MAIN-----------------------------------------------------------------------------------------
//##############################################################################################
//##############################################################################################
endmodule