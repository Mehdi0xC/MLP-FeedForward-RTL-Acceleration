// SYNTHESIZABLE MULTIPLIER FOR N BIT SIGNED MAGNITUDE WITH F BITS OF FRACTION
// CREATED BY MEHDI SAFAEE, WINTER 2018-2019
`include "config.svh"
module matrixMultiplier 
//##############################################################################################
//##############################################################################################
// PARAMETERs-----------------------------------------------------------------------------------
	#(
	parameter R = 3,
	parameter C = 4
	)
// INPUT AND OUTPUTS----------------------------------------------------------------------------
	(
	 input logic		[`N-1:0]	a[0:R-1],[`N-1:0] b[0:R-1][0:C-1],
	 output	logic		[`N-1:0]	c[0:R-1][0:C-1]
	 );
// VARIABLES -----------------------------------------------------------------------------------
	logic [`N-1:0] result[0:R-1][0:C-1];
	assign c = result;
// MODULES INSTANTIATIONS-----------------------------------------------------------------------
genvar i, j;
generate
	for (i=0; i<R; i=i+1) begin : loop_on_rows
	    for (j=0; j<C; j=j+1) begin : loop_on_columns
    multiplier multiplier_instance (
        .a(a[i]),
        .b(b[i][j]),
		.c(result[i][j])
    );
	end
	end
endgenerate
// INITIALIZATIONS------------------------------------------------------------------------------	
// MAIN-----------------------------------------------------------------------------------------
//##############################################################################################
//##############################################################################################
endmodule