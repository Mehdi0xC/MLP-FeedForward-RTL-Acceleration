// SYNTHESIZABLE ADDER FOR N BIT SIGNED MAGNITUDE WITH F BITS OF FRACTION
// CREATED BY MEHDI SAFAEE, WINTER 2018-2019
`include "config.svh"
module sigma32
//##############################################################################################
//##############################################################################################
// PARAMETERs-----------------------------------------------------------------------------------
// INPUT AND OUTPUTS----------------------------------------------------------------------------
    (
    input logic [`N-1:0] a[0:31][1],
    output logic [`N-1:0] c
    );
// MODULES INSTANTIATIONS-----------------------------------------------------------------------
    logic [`N-1:0] temp [0:1];
    logic [`N-1:0] result;
	sigma16 sigma16_0 
    (
		.a(a[0:15]), 
		.c(temp[0])
	);
    sigma16 sigma16_1
    (
		.a(a[16:31]), 
		.c(temp[1])
	);
	adder adder0
    (
		.a(temp[0]), 
		.b(temp[1]), 
		.c(result)
	);
// VARIABLES -----------------------------------------------------------------------------------
    assign c = result;
// INITIALIZATIONS------------------------------------------------------------------------------
// MAIN-----------------------------------------------------------------------------------------
//##############################################################################################
//##############################################################################################
endmodule