// MULTIPLYING PI AND NEPER NUMBER TOGETHER, WITH 32 BIT SIGNED MAGNITUDE REPRESENTATION AND 17 BIT OF FRACTIONS
// CREATED BY MEHDI SAFAEE, WINTER 2018-2019
`include "config.svh"
module mask_test;
//##############################################################################################
//##############################################################################################
// PARAMETERs-----------------------------------------------------------------------------------
    parameter R = 6;
	parameter C = 6;
// INPUT AND OUTPUTS----------------------------------------------------------------------------
// VARIABLES -----------------------------------------------------------------------------------
	 logic		[`N-1:0]	a[1][0:C-1];
     logic      [`N-1:0] b[0:R-1][0:C-1];
	 logic		[`N-1:0]	c[0:R-1][0:C-1];
     // MODULES INSTANTIATIONS-----------------------------------------------------------------------	
	mask #(.R(R), .C(C)) mask0 (
		.a(a), 
		.b(b), 
		.c(c)
	);
// INITIALIZATIONS------------------------------------------------------------------------------	
// MAIN-----------------------------------------------------------------------------------------
    always
    begin
        #100;
        a[0][0] = 32'h00ffffff;
        a[0][1] = 32'h00000000;		
        a[0][2] = 32'h00056fc2;		
        a[0][3] = 32'h00056fc2;		
        a[0][4] = 32'h00056fc2;		
        a[0][5] = 32'h00056fc2;		

        b[0][0] = 32'h0006487e;		
        b[0][1] = 32'h0006487e;		
        b[0][2] = 32'h0006487e;		
        b[0][3] = 32'h0006487e;		
        b[0][4] = 32'h0006487e;		
        b[0][5] = 32'h0006487e;		
        b[1][0] = 32'h0006487e;		
        b[1][1] = 32'h0006487e;		
        b[1][2] = 32'h0006487e;		
        b[1][3] = 32'h0006487e;		
        b[1][4] = 32'h0006487e;		
        b[1][5] = 32'h0006487e;		
        b[2][0] = 32'h0006487e;		
        b[2][1] = 32'h0006487e;		
        b[2][2] = 32'h0006487e;		
        b[2][3] = 32'h0006487e;		
        b[2][4] = 32'h0006487e;		
        b[2][5] = 32'h0006487e;		
        b[3][0] = 32'h0006487e;		
        b[3][1] = 32'h0006487e;		
        b[3][2] = 32'h0006487e;		
        b[3][3] = 32'h0006487e;		
        b[3][4] = 32'h0006487e;		
        b[3][5] = 32'h0006487e;		
        b[4][0] = 32'h0006487e;		
        b[4][1] = 32'h0006487e;		
        b[4][2] = 32'h0006487e;		
        b[4][3] = 32'h0006487e;		
        b[4][4] = 32'h0006487e;		
        b[4][5] = 32'h0006487e;		
        b[5][0] = 32'h0006487e;		
        b[5][1] = 32'h0006487e;		
        b[5][2] = 32'h0006487e;		
        b[5][3] = 32'h0006487e;		
        b[5][4] = 32'h0006487e;	
        b[5][5] = 32'h0006487e;		
	
    end
//##############################################################################################
//##############################################################################################
endmodule