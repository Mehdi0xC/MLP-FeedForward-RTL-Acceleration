// SYNTHESIZABLE ADDER FOR N BIT SIGNED MAGNITUDE WITH F BITS OF FRACTION
// CREATED BY MEHDI SAFAEE, WINTER 2018-2019
`include "config.svh"
module sigma7
//##############################################################################################
//##############################################################################################
// PARAMETERs-----------------------------------------------------------------------------------
// INPUT AND OUTPUTS----------------------------------------------------------------------------
    (
    input logic [`N-1:0] a[0:6][1],
    output logic [`N-1:0] c
    );
// MODULES INSTANTIATIONS-----------------------------------------------------------------------
    logic [`N-1:0] temp [0:4];
    logic [`N-1:0] result;

	adder adder0 
    (
		.a(a[0][0]), 
		.b(a[1][0]), 
		.c(temp[0])
	);
	adder adder1 
    (
		.a(a[2][0]), 
		.b(a[3][0]), 
		.c(temp[1])
	);
	adder adder2 
    (
		.a(a[4]), 
		.b(a[5]), 
		.c(temp[2])
	);
	adder adder3 
    (
		.a(a[6]), 
		.b(temp[2]), 
		.c(temp[4])
	);
	adder adder4 
    (
		.a(temp[0]), 
		.b(temp[1]), 
		.c(temp[3])
	);
	adder adder5 
    (
		.a(temp[3]), 
		.b(temp[4]), 
		.c(result)
	);
// VARIABLES -----------------------------------------------------------------------------------
    assign c = result;
// INITIALIZATIONS------------------------------------------------------------------------------
// MAIN-----------------------------------------------------------------------------------------
//##############################################################################################
//##############################################################################################
endmodule