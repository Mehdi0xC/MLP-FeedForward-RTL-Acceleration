`ifndef _config_svh_
`define _config_svh_
`define F 17
`define N 22
`define nNeurons 8
`define nActions 3
`define nStates 3
`define nSamples 100
`define nRewards 2
`endif
