// SYNTHESIZABLE ADDER FOR N BIT SIGNED MAGNITUDE WITH F BITS OF FRACTION
// CREATED BY MEHDI SAFAEE, WINTER 2018-2019
`include "config.svh"
module sigma4 
//##############################################################################################
//##############################################################################################
// PARAMETERs-----------------------------------------------------------------------------------
// INPUT AND OUTPUTS----------------------------------------------------------------------------
    (
    input logic [`N-1:0] a0, a1, a2, a3,
    output logic [`N-1:0] c
    );
// MODULES INSTANTIATIONS-----------------------------------------------------------------------
    logic [`N-1:0] temp [0:1];
    logic [`N-1:0] result;

	adder  adder0 
    (
		.a(a0), 
		.b(a1), 
		.c(temp[0])
	);
    adder  adder1 
    (
		.a(a2), 
		.b(a3), 
		.c(temp[1])
	);
	adder  adder2 
    (
		.a(temp[0]), 
		.b(temp[1]), 
		.c(result)
	);
// VARIABLES -----------------------------------------------------------------------------------
    assign c = result;
// INITIALIZATIONS------------------------------------------------------------------------------
// MAIN-----------------------------------------------------------------------------------------
//##############################################################################################
//##############################################################################################
endmodule