// ADDING PI AND NEPER NUMBER TOGETHER, WITH 32 BIT SIGNED MAGNITUDE REPRESENTATION AND 17 BIT OF FRACTIONS
// CREATED BY MEHDI SAFAEE, WINTER 2018-2019
`include "config.svh"
module sigma32_test;
//##############################################################################################
//##############################################################################################
// PARAMETERs-----------------------------------------------------------------------------------
// INPUT AND OUTPUTS----------------------------------------------------------------------------
// VARIABLES -----------------------------------------------------------------------------------
	logic [31:0] a[0:31][1];
	logic [31:0] c;
// MODULES INSTANTIATIONS-----------------------------------------------------------------------
	sigma32  sigma32_0 
    (
		.a(a), 
		.c(c)
	);
// INITIALIZATIONS------------------------------------------------------------------------------

// MAIN-----------------------------------------------------------------------------------------
    always
    begin
        #100;
        a[0][0] = 32'h0006487e;	
        a[1][0] = 32'h0006487e;		
        a[2][0] = 32'h0006487e;	
        a[3][0] = 32'h0006487e;	
        a[4][0] = 32'h0006487e;		
        a[5][0] = 32'h0006487e;	        	
        a[6][0] = 32'h0006487e;	        	
        a[7][0] = 32'h0006487e;	        	
        a[8][0] = 32'h0006487e;	        	
        a[9][0] = 32'h0006487e;	        	
        a[10][0] = 32'h0006487e;	        	
        a[11][0] = 32'h0006487e;	        	
        a[12][0] = 32'h0006487e;	        	
        a[13][0] = 32'h0006487e;	        	
        a[14][0] = 32'h0006487e;	        	
        a[15][0] = 32'h0006487e;	        	
        a[16][0] = 32'h0006487e;	        	
        a[17][0] = 32'h0006487e;	        	
        a[18][0] = 32'h0006487e;	        	
        a[19][0] = 32'h0006487e;	        	
        a[20][0] = 32'h0006487e;	        	
        a[21][0] = 32'h0006487e;	        	
        a[22][0] = 32'h0006487e;	        	
        a[23][0] = 32'h0006487e;	        	
        a[24][0] = 32'h0006487e;	        	
        a[25][0] = 32'h0006487e;	        	
        a[26][0] = 32'h0006487e;	        	
        a[27][0] = 32'h0006487e;	        	
        a[28][0] = 32'h0006487e;	        	
        a[29][0] = 32'h0006487e;	        	
        a[30][0] = 32'h0006487e;	        	
        a[31][0] = 32'h0006487e;	        	
    end
//##############################################################################################
//##############################################################################################
endmodule