// ADDING PI AND NEPER NUMBER TOGETHER, WITH 32 BIT SIGNED MAGNITUDE REPRESENTATION AND 17 BIT OF FRACTIONS
// CREATED BY MEHDI SAFAEE, WINTER 2018-2019
`include "config.svh"
module sigma_test;
//##############################################################################################
//##############################################################################################
// PARAMETERs-----------------------------------------------------------------------------------
// INPUT AND OUTPUTS----------------------------------------------------------------------------
// VARIABLES -----------------------------------------------------------------------------------
	logic [31:0] a[0:2][1];
	logic [31:0] c;
// MODULES INSTANTIATIONS-----------------------------------------------------------------------
	sigma3  sigma3_0 
    (
		.a(a), 
		.c(c)
	);
// INITIALIZATIONS------------------------------------------------------------------------------

// MAIN-----------------------------------------------------------------------------------------
    always
    begin
        #100;
        a[0][0] = 32'h0006487e;	
        a[1][0] = 32'h0006487e;		
        a[2][0] = 32'h0006487e;		
    end
//##############################################################################################
//##############################################################################################
endmodule